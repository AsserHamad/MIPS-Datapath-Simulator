module main()
